module vga_controller

endmodule 