
`include "uart_tx.v"
`include "uart_rx.v"
`include "vga_controller"

module main(
    input;
    output;
    );
    
    //Check signal from UART
    
    //check sinal of putput
endmodule
