
`timescale 1ns/10ps

`include "vga_controller.v"

module vga_tb();
    
endmodule