
`include "uart_tx.v"
`include "uart_rx.v"
`include "vga_controller"

module main
endmodule
